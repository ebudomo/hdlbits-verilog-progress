module wire_simple( 
	input in, 
	output out 
);
    
	assign out = in;

endmodule 