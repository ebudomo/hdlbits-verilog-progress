module circuit1(
	input a,
	input b,
	output q
);

endmodule
