module circuit1(
	input a,
	input b,
	output q
);
	// waveform displays circuit that implements q = a & b
	assign q = a & b;

endmodule
