module m2014_q4h(
	input in,
	output out
);
	// implement a simple wire connecting input and output ports
	assign out = in;
	
endmodule
