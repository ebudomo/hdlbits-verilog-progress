module m2014_q4i(
	output out
);
	// implement an output port set to ground
	assign out = 1'b0;

endmodule
