library verilog;
use verilog.vl_types.all;
entity clock is
end clock;
