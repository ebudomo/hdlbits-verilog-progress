module dut ( input clk, output q ) ;
	// provided module
	assign q = clk;
	
endmodule
